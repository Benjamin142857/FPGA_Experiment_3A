-------------------------------------------------------------------------------
-- Title         : rom lookup table
-- Project       : umts_interleaver
-------------------------------------------------------------------------------
-- File          : $Workfile:   aukui_prime_rom_e.vhd  $
-- Revision      : $Revision: #1 $
-- Author        : Volker Mauer
-- Checked in by : $Author: zpan $
-- Last modified : $Date: 2009/06/19 $
-------------------------------------------------------------------------------
-- Description :
--
-- ROM containing prime numbers and primitive roots
--
-- Copyright 2000 (c) Altera Corporation
-- All rights reserved
--
-------------------------------------------------------------------------------
-- Modification history :
-- $Log: $
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library auk_dspip_ctc_umts_lib;
use auk_dspip_ctc_umts_lib.auk_dspip_ctc_umts_lib_pkg.all;

entity auk_dspip_ctc_umtsitlv_prime_rom is

    port (
        prime_index : in unsigned(6 downto 0);

        prime : out unsigned(8 downto 0);
        g0    : out unsigned(4 downto 0);
-- gcd : out vec_of_vec(19 downto 0, 5 downto 0);
-- gcd : out gcd_vec;

        gcd_index : in  unsigned(4 downto 0);
        gcd       : out unsigned(7 downto 0);

        reset  : in std_logic;
        enable : in std_logic;
        clk    : in std_logic
        );

end auk_dspip_ctc_umtsitlv_prime_rom;



architecture beh of auk_dspip_ctc_umtsitlv_prime_rom is

    type gcd_vec is array (19 downto 0) of unsigned(7 downto 0);

    signal rd_addr_int : integer;
    signal primevec    : std_logic_vector(45 downto 12);
    signal gcd_int     : gcd_vec;
    signal primeval    : unsigned(8 downto 0);
    signal g0val       : unsigned(4 downto 0);
    signal gcdval      : unsigned(139 downto 0);

begin  -- beh

    rd_addr_int <= to_integer(prime_index);

    gcd <= gcd_int(to_integer(gcd_index));


    prime_lookup : process (rd_addr_int)

    begin  -- process lookup
        case rd_addr_int is
            when 0      => primeval <= "000000111";  -- dummy line
            when 1      => primeval <= "000000111";  -- dummy line
            when 2      => primeval <= "000000111";
            when 3      => primeval <= "000001011";
            when 4      => primeval <= "000001101";
            when 5      => primeval <= "000010001";
            when 6      => primeval <= "000010011";
            when 7      => primeval <= "000010111";
            when 8      => primeval <= "000011101";
            when 9      => primeval <= "000011111";
            when 10     => primeval <= "000100101";
            when 11     => primeval <= "000101001";
            when 12     => primeval <= "000101011";
            when 13     => primeval <= "000101111";
            when 14     => primeval <= "000110101";
            when 15     => primeval <= "000111011";
            when 16     => primeval <= "000111101";
            when 17     => primeval <= "001000011";
            when 18     => primeval <= "001000111";
            when 19     => primeval <= "001001001";
            when 20     => primeval <= "001001111";
            when 21     => primeval <= "001010011";  -- 97
            when 22     => primeval <= "001011001";
            when 23     => primeval <= "001100001";
            when 24     => primeval <= "001100101";
            when 25     => primeval <= "001100111";
            when 26     => primeval <= "001101011";
            when 27     => primeval <= "001101101";
            when 28     => primeval <= "001110001";
            when 29     => primeval <= "001111111";
            when 30     => primeval <= "010000011";
            when 31     => primeval <= "010001001";
            when 32     => primeval <= "010001011";
            when 33     => primeval <= "010010101";
            when 34     => primeval <= "010010111";
            when 35     => primeval <= "010011101";
            when 36     => primeval <= "010100011";
            when 37     => primeval <= "010100111";
            when 38     => primeval <= "010101101";
            when 39     => primeval <= "010110011";
            when 40     => primeval <= "010110101";
            when 41     => primeval <= "010111111";
            when 42     => primeval <= "011000001";
            when 43     => primeval <= "011000101";  -- 211
            when 44     => primeval <= "011000111";
            when 45     => primeval <= "011010011";
            when 46     => primeval <= "011011111";
            when 47     => primeval <= "011100011";
            when 48     => primeval <= "011100101";
            when 49     => primeval <= "011101001";
            when 50     => primeval <= "011101111";
            when 51     => primeval <= "011110001";
            when 52     => primeval <= "011111011";
            when 53     => primeval <= "100000001";
            when others => primeval <= "---------";  -- dummy line
        end case;
    end process prime_lookup;

    gcd_lookup : process (rd_addr_int)

    begin  -- process lookup
        case rd_addr_int is
            when 0      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- dummy line
            when 1      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- dummy line
            when 2      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 7
            when 3      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 11
            when 4      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 13
            when 5      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 17
            when 6      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 19
            when 7      => gcdval <= "00000010000111000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 23
            when 8      => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 29
            when 9      => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 31
            when 10     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 37
            when 11     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 41
            when 12     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 43
            when 13     => gcdval <= "00000010000111000101100011010010001001001100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 47
            when 14     => gcdval <= "00000010000111000101100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 53
            when 15     => gcdval <= "00000010000111000101100011010010001001001100101110011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 59
            when 16     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 61
            when 17     => gcdval <= "00000010000111000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 67
            when 18     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 71
            when 19     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 73
            when 20     => gcdval <= "00000010000111000101100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 79
            when 21     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101011010111101101010111011011110110000111000111100100110011111010011";  -- 83
            when 22     => gcdval <= "00000010000111000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 89
            when 23     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 97
            when 24     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 101
            when 25     => gcdval <= "00000010000111000101100011010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 103
            when 26     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110111011011110110000111000111100100110011111010011";  -- 107
            when 27     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 109
            when 28     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 113
            when 29     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 127
            when 30     => gcdval <= "00000010000111000101100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 131
            when 31     => gcdval <= "00000010000111000101100011010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 137
            when 32     => gcdval <= "00000010000111000101100011010010001001001100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 139
            when 33     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 149
            when 34     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 151
            when 35     => gcdval <= "00000010000111000101100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 157
            when 36     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 163
            when 37     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 167
            when 38     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010111101101010111011011110110000111000111100100110011111010011";  -- 173
            when 39     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 179
            when 40     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 181
            when 41     => gcdval <= "00000010000111000101100011010010001001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 191
            when 42     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 193
            when 43     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 197
            when 44     => gcdval <= "00000010000111000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 199
            when 45     => gcdval <= "00000010001011000110100100010010011001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 211
            when 46     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 223
            when 47     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 227
            when 48     => gcdval <= "00000010000111000101100011010010001001011100111010011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 229
            when 49     => gcdval <= "00000010000111000101100011010010001001001100101110011111010010101010010101011010111101101010111011011110110000111000111100100110011111010011";  -- 233
            when 50     => gcdval <= "00000010001011000110100100110010111001110100111110100101010100101010110101111011010101110110111101100001110001111001001100111110100111011001";  -- 239
            when 51     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 241
            when 52     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 251
            when 53     => gcdval <= "00000010000111000101100011010010001001001100101110011101001111101001010101001010101101011110110101011101101111011000011100011110010011001111";  -- 257
            when others => gcdval <= "--------------------------------------------------------------------------------------------------------------------------------------------";  -- dummy line
--        when  0 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- dummy line
--        when  1 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- dummy line
--        when  2 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 7
--        when  3 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 11
--        when  4 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 13
--        when  5 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 17
--        when  6 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 19
--        when  7 => gcdval <= "1,7,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 23
--        when  8 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 29
--        when  9 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 31
--        when 10 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 37
--        when 11 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 41
--        when 12 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 43
--        when 13 => gcdval <= "1,7,11,13,17,19,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 47
--        when 14 => gcdval <= "1,7,11,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 53
--        when 15 => gcdval <= "1,7,11,13,17,19,23,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 59
--        when 16 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 61
--        when 17 => gcdval <= "1,7,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 67
--        when 18 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 71
--        when 19 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 73
--        when 20 => gcdval <= "1,7,11,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 79
--        when 21 => gcdval <= "1,7,11,13,17,19,23,29,31,37,43,47,53,59,61,67,71,73,79,83,89";  -- 83
--        when 22 => gcdval <= "1,7,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 89
--        when 23 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 97
--        when 24 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 101
--        when 25 => gcdval <= "1,7,11,13,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 103
--        when 26 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,59,61,67,71,73,79,83,89";  -- 107
--        when 27 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 109
--        when 28 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 113
--        when 29 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 127
--        when 30 => gcdval <= "1,7,11,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 131
--        when 31 => gcdval <= "1,7,11,13,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 137
--        when 32 => gcdval <= "1,7,11,13,17,19,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 139
--        when 33 => gcdval <= "1,7,11,13,17,19,23,29,31,41,43,47,53,59,61,67,71,73,79,83,89";  -- 149
--        when 34 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 151
--        when 35 => gcdval <= "1,7,11,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 157
--        when 36 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 163
--        when 37 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,89";  -- 167
--        when 38 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,47,53,59,61,67,71,73,79,83,89";  -- 173
--        when 39 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 179
--        when 40 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 181
--        when 41 => gcdval <= "1,7,11,13,17,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 191
--        when 42 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 193
--        when 43 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 197
--        when 44 => gcdval <= "1,7,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 199
--        when 45 => gcdval <= "1,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 211
--        when 46 => gcdval <= "1,7,11,13,17,19,23,29,31,41,43,47,53,59,61,67,71,73,79,83,89";  -- 223
--        when 47 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 227
--        when 48 => gcdval <= "1,7,11,13,17,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 229
--        when 49 => gcdval <= "1,7,11,13,17,19,23,31,37,41,43,47,53,59,61,67,71,73,79,83,89";  -- 233
--        when 50 => gcdval <= "1,11,13,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83,89,97";  -- 239
--        when 51 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 241
--        when 52 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 251
--        when 53 => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- 257
--    when others => gcdval <= "1,7,11,13,17,19,23,29,31,37,41,43,47,53,59,61,67,71,73,79,83";  -- dummy line
        end case;
    end process gcd_lookup;

    g0_lookup : process (rd_addr_int)

    begin  -- process lookup
        case rd_addr_int is
            when 0      => g0val <= "00011";  -- dummy line
            when 1      => g0val <= "00011";  -- dummy line
            when 2      => g0val <= "00011";
            when 3      => g0val <= "00010";
            when 4      => g0val <= "00010";
            when 5      => g0val <= "00011";
            when 6      => g0val <= "00010";
            when 7      => g0val <= "00101";
            when 8      => g0val <= "00010";
            when 9      => g0val <= "00011";
            when 10     => g0val <= "00010";
            when 11     => g0val <= "00110";
            when 12     => g0val <= "00011";
            when 13     => g0val <= "00101";
            when 14     => g0val <= "00010";
            when 15     => g0val <= "00010";
            when 16     => g0val <= "00010";
            when 17     => g0val <= "00010";
            when 18     => g0val <= "00111";
            when 19     => g0val <= "00101";
            when 20     => g0val <= "00011";
            when 21     => g0val <= "00010";  -- 97
            when 22     => g0val <= "00011";
            when 23     => g0val <= "00101";
            when 24     => g0val <= "00010";
            when 25     => g0val <= "00101";
            when 26     => g0val <= "00010";
            when 27     => g0val <= "00110";
            when 28     => g0val <= "00011";
            when 29     => g0val <= "00011";
            when 30     => g0val <= "00010";
            when 31     => g0val <= "00011";
            when 32     => g0val <= "00010";
            when 33     => g0val <= "00010";
            when 34     => g0val <= "00110";
            when 35     => g0val <= "00101";
            when 36     => g0val <= "00010";
            when 37     => g0val <= "00101";
            when 38     => g0val <= "00010";
            when 39     => g0val <= "00010";
            when 40     => g0val <= "00010";
            when 41     => g0val <= "10011";
            when 42     => g0val <= "00101";
            when 43     => g0val <= "00010";  -- 211
            when 44     => g0val <= "00011";
            when 45     => g0val <= "00010";
            when 46     => g0val <= "00011";
            when 47     => g0val <= "00010";
            when 48     => g0val <= "00110";
            when 49     => g0val <= "00011";
            when 50     => g0val <= "00111";
            when 51     => g0val <= "00111";
            when 52     => g0val <= "00110";
            when 53     => g0val <= "00011";
            when others => g0val <= "-----";  -- dummy line
        end case;
    end process g0_lookup;


    -- purpose: <description>
    out_signals : process (clk, reset)
        
    begin  -- process out_signals
        -- activities triggered by asynchronous reset (active high)
        if reset = '1' then
            prime <= (others => '0');
            g0 <= (others => '0');
            reset_loop : for i in 0 to 19 loop
                gcd_int(i) <= (others => '0');
            end loop reset_loop;
            -- activities triggered by rising edge of clock
        elsif clk'event and clk = '1' then
            if enable = '1' then
                
                if rd_addr_int < 2 then
                    prime <= to_unsigned(0,9);
                else
                    prime <= primeval;
--		    prime <= ('0' & unsigned(primevec(45 downto 39))) & '0' + to_unsigned(17, 9);
--		    prime <= ('0' & unsigned(primevec(45 downto 39))) & '1' + to_unsigned(16, 9);  -- should synthesize better
                end if;

                g0 <= g0val;

                out_loop : for i in 0 to 19 loop
                    gcd_int(i) <= '0' & gcdval((19-i)*7+6 downto (19-i)*7+0);
--		    gcd_int(i) <= '0' & gcdval(i*7+6 downto i*7+0);
                end loop out_loop;
                
            end if;
            
        end if;
    end process out_signals;
end beh;
