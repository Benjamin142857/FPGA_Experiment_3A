-- megafunction wizard: %ALTMULT_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTMULT_ADD 

-- ============================================================
-- File Name: four_mult_add.vhd
-- Megafunction Name(s):
-- 			ALTMULT_ADD
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--Copyright (C) 1991-2003 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY four_mult_add IS
	PORT
	(
		clock0		: IN STD_LOGIC  := '1';
		dataa_0		: IN STD_LOGIC_VECTOR (15 DOWNTO 0) :=  (OTHERS => '0');
		aclr3		: IN STD_LOGIC  := '0';
		datab_0		: IN STD_LOGIC_VECTOR (13 DOWNTO 0) :=  (OTHERS => '0');
		datab_1		: IN STD_LOGIC_VECTOR (13 DOWNTO 0) :=  (OTHERS => '0');
		datab_2		: IN STD_LOGIC_VECTOR (13 DOWNTO 0) :=  (OTHERS => '0');
		datab_3		: IN STD_LOGIC_VECTOR (13 DOWNTO 0) :=  (OTHERS => '0');
		shiftouta		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END four_mult_add;


ARCHITECTURE SYN OF four_mult_add IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire2_bv	: BIT_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (63 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (55 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (13 DOWNTO 0);



	COMPONENT altmult_add
	GENERIC (
		input_register_b2		: STRING;
		input_register_a1		: STRING;
		multiplier_register0		: STRING;
		signed_pipeline_aclr_b		: STRING;
		input_register_b3		: STRING;
		input_register_a2		: STRING;
		multiplier_register1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		input_register_a3		: STRING;
		multiplier_register2		: STRING;
		signed_aclr_a		: STRING;
		signed_register_a		: STRING;
		number_of_multipliers		: NATURAL;
		multiplier_register3		: STRING;
		multiplier_aclr0		: STRING;
		addnsub_multiplier_pipeline_aclr3		: STRING;
		signed_aclr_b		: STRING;
		signed_register_b		: STRING;
		lpm_type		: STRING;
		multiplier_aclr1		: STRING;
		input_aclr_b0		: STRING;
		output_register		: STRING;
		representation_a		: STRING;
		signed_pipeline_register_a		: STRING;
		width_result		: NATURAL;
		input_source_b0		: STRING;
		multiplier_aclr2		: STRING;
		input_aclr_b1		: STRING;
		input_aclr_a0		: STRING;
		multiplier3_direction		: STRING;
		addnsub_multiplier_register1		: STRING;
		representation_b		: STRING;
		signed_pipeline_register_b		: STRING;
		input_source_b1		: STRING;
		input_source_a0		: STRING;
		multiplier_aclr3		: STRING;
		input_aclr_b2		: STRING;
		input_aclr_a1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_source_b2		: STRING;
		input_source_a1		: STRING;
		input_aclr_b3		: STRING;
		input_aclr_a2		: STRING;
		addnsub_multiplier_register3		: STRING;
		addnsub_multiplier_aclr1		: STRING;
		output_aclr		: STRING;
		input_source_b3		: STRING;
		input_source_a2		: STRING;
		input_aclr_a3		: STRING;
		input_source_a3		: STRING;
		addnsub_multiplier_aclr3		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		width_a		: NATURAL;
		input_register_b0		: STRING;
		width_b		: NATURAL;
		input_register_b1		: STRING;
		input_register_a0		: STRING;
		addnsub_multiplier_pipeline_register3		: STRING;
		multiplier1_direction		: STRING;
		signed_pipeline_aclr_a		: STRING
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (55 DOWNTO 0);
			scanouta	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire2_bv(15 DOWNTO 0) <= "0000000000000000";
	sub_wire2    <= To_stdlogicvector(sub_wire2_bv);
	shiftouta    <= sub_wire0(15 DOWNTO 0);
	result    <= sub_wire1(31 DOWNTO 0);
	sub_wire4    <= dataa_0(15 DOWNTO 0);
	sub_wire3    <= sub_wire2(15 DOWNTO 0) & sub_wire2(15 DOWNTO 0) & sub_wire2(15 DOWNTO 0) & sub_wire4(15 DOWNTO 0);
	sub_wire5    <= datab_1(13 DOWNTO 0);
	sub_wire7    <= datab_0(13 DOWNTO 0);
	sub_wire8    <= datab_2(13 DOWNTO 0);
	sub_wire9    <= datab_3(13 DOWNTO 0);
	sub_wire6    <= sub_wire9(13 DOWNTO 0) & sub_wire8(13 DOWNTO 0) & sub_wire5(13 DOWNTO 0) & sub_wire7(13 DOWNTO 0);

	ALTMULT_ADD_component : altmult_add
	GENERIC MAP (
		input_register_b2 => "CLOCK0",
		input_register_a1 => "CLOCK0",
		multiplier_register0 => "CLOCK0",
		signed_pipeline_aclr_b => "ACLR3",
		input_register_b3 => "CLOCK0",
		input_register_a2 => "CLOCK0",
		multiplier_register1 => "CLOCK0",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		input_register_a3 => "CLOCK0",
		multiplier_register2 => "CLOCK0",
		signed_aclr_a => "ACLR3",
		signed_register_a => "CLOCK0",
		number_of_multipliers => 4,
		multiplier_register3 => "CLOCK0",
		multiplier_aclr0 => "ACLR3",
		addnsub_multiplier_pipeline_aclr3 => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_register_b => "CLOCK0",
		lpm_type => "altmult_add",
		multiplier_aclr1 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		output_register => "CLOCK0",
		representation_a => "SIGNED",
		signed_pipeline_register_a => "CLOCK0",
		width_result => 32,
		input_source_b0 => "DATAB",
		multiplier_aclr2 => "ACLR3",
		input_aclr_b1 => "ACLR3",
		input_aclr_a0 => "ACLR3",
		multiplier3_direction => "ADD",
		addnsub_multiplier_register1 => "CLOCK0",
		representation_b => "SIGNED",
		signed_pipeline_register_b => "CLOCK0",
		input_source_b1 => "DATAB",
		input_source_a0 => "SCANA",
		multiplier_aclr3 => "ACLR3",
		input_aclr_b2 => "ACLR3",
		input_aclr_a1 => "ACLR3",
		dedicated_multiplier_circuitry => "YES",
		input_source_b2 => "DATAB",
		input_source_a1 => "SCANA",
		input_aclr_b3 => "ACLR3",
		input_aclr_a2 => "ACLR3",
		addnsub_multiplier_register3 => "CLOCK0",
		addnsub_multiplier_aclr1 => "ACLR3",
		output_aclr => "ACLR3",
		input_source_b3 => "DATAB",
		input_source_a2 => "SCANA",
		input_aclr_a3 => "ACLR3",
		input_source_a3 => "SCANA",
		addnsub_multiplier_aclr3 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		width_a => 16,
		input_register_b0 => "CLOCK0",
		width_b => 14,
		input_register_b1 => "CLOCK0",
		input_register_a0 => "CLOCK0",
		addnsub_multiplier_pipeline_register3 => "CLOCK0",
		multiplier1_direction => "ADD",
		signed_pipeline_aclr_a => "ACLR3"
	)
	PORT MAP (
		dataa => sub_wire3,
		datab => sub_wire6,
		clock0 => clock0,
		aclr3 => aclr3,
		scanouta => sub_wire0,
		result => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: SRCA0 STRING "Shiftin input"
-- Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNA STRING "Signed"
-- Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: MULT_REGOUT0 STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB STRING "Signed"
-- Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: SAME_CONFIG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGB0 STRING "1"
-- Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGA0 STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED STRING "1"
-- Retrieval info: PRIVATE: RTS_WIDTH STRING "32"
-- Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: IMPL_STYLE_LCELL STRING "0"
-- Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: NUM_MULT STRING "4"
-- Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: SCANOUTA STRING "1"
-- Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: REG_OUT STRING "1"
-- Retrieval info: PRIVATE: SCANOUTB STRING "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT STRING "0"
-- Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADD_ENABLE STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ALL_REG_ACLR STRING "1"
-- Retrieval info: PRIVATE: WIDTHA STRING "16"
-- Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_REG STRING "1"
-- Retrieval info: PRIVATE: WIDTHB STRING "14"
-- Retrieval info: PRIVATE: SIGNB_REG STRING "1"
-- Retrieval info: PRIVATE: OP1 STRING "Add"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: OP3 STRING "Add"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INPUT_REGISTER_B2 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_B STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B3 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A2 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A3 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER2 STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_ACLR_A STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "4"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER3 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR0 STRING "ACLR3"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR3 STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_ACLR_B STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_B0 STRING "ACLR3"
-- Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR2 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_B1 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_A0 STRING "ACLR3"
-- Retrieval info: CONSTANT: MULTIPLIER3_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "SCANA"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR3 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_B2 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_A1 STRING "ACLR3"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B2 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "SCANA"
-- Retrieval info: CONSTANT: INPUT_ACLR_B3 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_A2 STRING "ACLR3"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER3 STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: OUTPUT_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B3 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A2 STRING "SCANA"
-- Retrieval info: CONSTANT: INPUT_ACLR_A3 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A3 STRING "SCANA"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR3 STRING "ACLR3"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "14"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER3 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_A STRING "ACLR3"
-- Retrieval info: USED_PORT: shiftouta 0 0 16 0 OUTPUT GND "shiftouta[15..0]"
-- Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
-- Retrieval info: USED_PORT: dataa_0 0 0 16 0 INPUT GND "dataa_0[15..0]"
-- Retrieval info: USED_PORT: aclr3 0 0 0 0 INPUT GND "aclr3"
-- Retrieval info: USED_PORT: datab_0 0 0 14 0 INPUT GND "datab_0[13..0]"
-- Retrieval info: USED_PORT: datab_1 0 0 14 0 INPUT GND "datab_1[13..0]"
-- Retrieval info: USED_PORT: datab_2 0 0 14 0 INPUT GND "datab_2[13..0]"
-- Retrieval info: USED_PORT: datab_3 0 0 14 0 INPUT GND "datab_3[13..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT GND "result[31..0]"
-- Retrieval info: CONNECT: @datab 0 0 14 14 datab_1 0 0 14 0
-- Retrieval info: CONNECT: @datab 0 0 14 28 datab_2 0 0 14 0
-- Retrieval info: CONNECT: @datab 0 0 14 42 datab_3 0 0 14 0
-- Retrieval info: CONNECT: @aclr3 0 0 0 0 aclr3 0 0 0 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 16 48 GND 0 0 16 0
-- Retrieval info: CONNECT: @dataa 0 0 16 32 GND 0 0 16 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: CONNECT: @dataa 0 0 16 0 dataa_0 0 0 16 0
-- Retrieval info: CONNECT: @dataa 0 0 16 16 GND 0 0 16 0
-- Retrieval info: CONNECT: shiftouta 0 0 16 0 @scanouta 0 0 16 0
-- Retrieval info: CONNECT: @datab 0 0 14 0 datab_0 0 0 14 0
